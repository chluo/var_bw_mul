/* ======================================================================
 *
 * Half Adder
 *
 * ======================================================================
 * Basic Inforation 
 * ----------------------------------------------------------------------
 * Author           |  Chunheng Luo
 * ----------------------------------------------------------------------
 * Email Address    |  Chunheng.Luo@utexas.edu
 * ----------------------------------------------------------------------
 * Data of Creation |  04-16-2017
 * ----------------------------------------------------------------------
 * Description      |  Half adder
 * =================================================================== */

 module half_adder 
 ( 
   input   a  ,
   input   b  ,
   output  s  ,
   output  co  
 ) ;

   assign { co , s } = a + b ;

 endmodule 

