/* ======================================================================
 *
 * Full Adder
 *
 * ======================================================================
 * Basic Inforation 
 * ----------------------------------------------------------------------
 * Author           |  Chunheng Luo
 * ----------------------------------------------------------------------
 * Email Address    |  Chunheng.Luo@utexas.edu
 * ----------------------------------------------------------------------
 * Data of Creation |  04-16-2017
 * ----------------------------------------------------------------------
 * Description      |  Full adder
 * =================================================================== */

 module full_adder 
 ( 
   input   a  ,
   input   b  ,
   input   ci ,
   output  s  ,
   output  co  
 ) ;

   assign { co , s } = a + b + ci ;

 endmodule 
