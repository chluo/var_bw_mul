/* ======================================================================
 *
 * Fixed Bit-width 16-bit Array Multiplier (array_fix_bw_mul)
 *
 * ======================================================================
 * Basic Inforation 
 * ----------------------------------------------------------------------
 * Author           |  Wei Ye
 * ----------------------------------------------------------------------
 * Email Address    |  weiye@utexas.edu
 * ----------------------------------------------------------------------
 * Data of Creation |  04-13-2017
 * ----------------------------------------------------------------------
 * Description      |  16-bit array multiplier. 
 * =================================================================== */

 module array_var_bw_mul
 (
   input                 para_mode    , 
   input    [ 15 : 0 ]   a            , // Operand A 
   input    [ 15 : 0 ]   b            , // Operand B 
   output   [ 31 : 0 ]   p              // Product 
 ) ; 

   //
   // Internal signals 
   //
   // The stage outputs are aligned
   // The first matrix coming out from the AND gates (16 rows)
   wire     [ 15 : 0 ]   b_00_a  ; // Row  0
   wire     [ 15 : 0 ]   b_01_a  ; // Row  1
   wire     [ 15 : 0 ]   b_02_a  ; // Row  2
   wire     [ 15 : 0 ]   b_03_a  ; // Row  3
   wire     [ 15 : 0 ]   b_04_a  ; // Row  4
   wire     [ 15 : 0 ]   b_05_a  ; // Row  5
   wire     [ 15 : 0 ]   b_06_a  ; // Row  6
   wire     [ 15 : 0 ]   b_07_a  ; // Row  7
   wire     [ 15 : 0 ]   b_08_a  ; // Row  8
   wire     [ 15 : 0 ]   b_09_a  ; // Row  9
   wire     [ 15 : 0 ]   b_10_a  ; // Row 10
   wire     [ 15 : 0 ]   b_11_a  ; // Row 11
   wire     [ 15 : 0 ]   b_12_a  ; // Row 12
   wire     [ 15 : 0 ]   b_13_a  ; // Row 13
   wire     [ 15 : 0 ]   b_14_a  ; // Row 14
   wire     [ 15 : 0 ]   b_15_a  ; // Row 15

   //
   // AND's
   // 
   assign b_00_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  0 ] } } ;  
   assign b_01_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  1 ] } } ;  
   assign b_02_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  2 ] } } ;  
   assign b_03_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  3 ] } } ;  
   assign b_04_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  4 ] } } ;  
   assign b_05_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  5 ] } } ;  
   assign b_06_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  6 ] } } ;  
   assign b_07_a = ( para_mode ? { { 8 { 1'b0 } } , a [  7 : 0 ] } : a ) & { 16 { b [  7 ] } } ;  
   assign b_08_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [  8 ] } } ;  
   assign b_09_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [  9 ] } } ;  
   assign b_10_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 10 ] } } ;  
   assign b_11_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 11 ] } } ;  
   assign b_12_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 12 ] } } ;  
   assign b_13_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 13 ] } } ;  
   assign b_14_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 14 ] } } ;  
   assign b_15_a = ( para_mode ? { a [ 15 : 8 ] , { 8 { 1'b0 } } } : a ) & { 16 { b [ 15 ] } } ;  
 
    assign p [ 0 ] = b_00_a [ 0 ] ;

    //
    // Row 0
    //
    wire [ 1 : 0 ] fa_00_01 =                 b_01_a [  0 ] + b_00_a [  1 ] ;
    wire [ 1 : 0 ] fa_00_02 = b_02_a [  0 ] + b_01_a [  1 ] + b_00_a [  2 ] ;
    wire [ 1 : 0 ] fa_00_03 = b_02_a [  1 ] + b_01_a [  2 ] + b_00_a [  3 ] ;
    wire [ 1 : 0 ] fa_00_04 = b_02_a [  2 ] + b_01_a [  3 ] + b_00_a [  4 ] ;
    wire [ 1 : 0 ] fa_00_05 = b_02_a [  3 ] + b_01_a [  4 ] + b_00_a [  5 ] ;
    wire [ 1 : 0 ] fa_00_06 = b_02_a [  4 ] + b_01_a [  5 ] + b_00_a [  6 ] ;
    wire [ 1 : 0 ] fa_00_07 = b_02_a [  5 ] + b_01_a [  6 ] + b_00_a [  7 ] ;
    wire [ 1 : 0 ] fa_00_08 = b_02_a [  6 ] + b_01_a [  7 ] + b_00_a [  8 ] ;
    wire [ 1 : 0 ] fa_00_09 = b_02_a [  7 ] + b_01_a [  8 ] + b_00_a [  9 ] ;
    wire [ 1 : 0 ] fa_00_10 = b_02_a [  8 ] + b_01_a [  9 ] + b_00_a [ 10 ] ;
    wire [ 1 : 0 ] fa_00_11 = b_02_a [  9 ] + b_01_a [ 10 ] + b_00_a [ 11 ] ;
    wire [ 1 : 0 ] fa_00_12 = b_02_a [ 10 ] + b_01_a [ 11 ] + b_00_a [ 12 ] ;
    wire [ 1 : 0 ] fa_00_13 = b_02_a [ 11 ] + b_01_a [ 12 ] + b_00_a [ 13 ] ;
    wire [ 1 : 0 ] fa_00_14 = b_02_a [ 12 ] + b_01_a [ 13 ] + b_00_a [ 14 ] ;
    wire [ 1 : 0 ] fa_00_15 = b_02_a [ 13 ] + b_01_a [ 14 ] + b_00_a [ 15 ] ;

    assign p [ 1 ] = fa_00_01 [ 0 ] ;


   //
   // Row 1
   //
   wire [ 1 : 0 ] fa_01_02 = fa_00_01 [ 1 ] + fa_00_02 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_01_03 = fa_00_02 [ 1 ] + fa_00_03 [ 0 ] + b_03_a [  0 ] ;
   wire [ 1 : 0 ] fa_01_04 = fa_00_03 [ 1 ] + fa_00_04 [ 0 ] + b_03_a [  1 ] ;
   wire [ 1 : 0 ] fa_01_05 = fa_00_04 [ 1 ] + fa_00_05 [ 0 ] + b_03_a [  2 ] ;
   wire [ 1 : 0 ] fa_01_06 = fa_00_05 [ 1 ] + fa_00_06 [ 0 ] + b_03_a [  3 ] ;
   wire [ 1 : 0 ] fa_01_07 = fa_00_06 [ 1 ] + fa_00_07 [ 0 ] + b_03_a [  4 ] ;
   wire [ 1 : 0 ] fa_01_08 = fa_00_07 [ 1 ] + fa_00_08 [ 0 ] + b_03_a [  5 ] ;
   wire [ 1 : 0 ] fa_01_09 = fa_00_08 [ 1 ] + fa_00_09 [ 0 ] + b_03_a [  6 ] ;
   wire [ 1 : 0 ] fa_01_10 = fa_00_09 [ 1 ] + fa_00_10 [ 0 ] + b_03_a [  7 ] ;
   wire [ 1 : 0 ] fa_01_11 = fa_00_10 [ 1 ] + fa_00_11 [ 0 ] + b_03_a [  8 ] ;
   wire [ 1 : 0 ] fa_01_12 = fa_00_11 [ 1 ] + fa_00_12 [ 0 ] + b_03_a [  9 ] ;
   wire [ 1 : 0 ] fa_01_13 = fa_00_12 [ 1 ] + fa_00_13 [ 0 ] + b_03_a [ 10 ] ;
   wire [ 1 : 0 ] fa_01_14 = fa_00_13 [ 1 ] + fa_00_14 [ 0 ] + b_03_a [ 11 ] ;
   wire [ 1 : 0 ] fa_01_15 = fa_00_14 [ 1 ] + fa_00_15 [ 0 ] + b_03_a [ 12 ] ;
   wire [ 1 : 0 ] fa_01_16 = fa_00_15 [ 1 ] +  b_01_a [ 15 ] + b_02_a [ 14 ] ;
   
   assign p [ 2 ] = fa_01_02 [ 0 ] ;


   //
   // Row 2
   //
   wire [ 1 : 0 ] fa_02_03 = fa_01_02 [ 1 ] + fa_01_03 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_02_04 = fa_01_03 [ 1 ] + fa_01_04 [ 0 ] + b_04_a [  0 ] ;
   wire [ 1 : 0 ] fa_02_05 = fa_01_04 [ 1 ] + fa_01_05 [ 0 ] + b_04_a [  1 ] ;
   wire [ 1 : 0 ] fa_02_06 = fa_01_05 [ 1 ] + fa_01_06 [ 0 ] + b_04_a [  2 ] ;
   wire [ 1 : 0 ] fa_02_07 = fa_01_06 [ 1 ] + fa_01_07 [ 0 ] + b_04_a [  3 ] ;
   wire [ 1 : 0 ] fa_02_08 = fa_01_07 [ 1 ] + fa_01_08 [ 0 ] + b_04_a [  4 ] ;
   wire [ 1 : 0 ] fa_02_09 = fa_01_08 [ 1 ] + fa_01_09 [ 0 ] + b_04_a [  5 ] ;
   wire [ 1 : 0 ] fa_02_10 = fa_01_09 [ 1 ] + fa_01_10 [ 0 ] + b_04_a [  6 ] ;
   wire [ 1 : 0 ] fa_02_11 = fa_01_10 [ 1 ] + fa_01_11 [ 0 ] + b_04_a [  7 ] ;
   wire [ 1 : 0 ] fa_02_12 = fa_01_11 [ 1 ] + fa_01_12 [ 0 ] + b_04_a [  8 ] ;
   wire [ 1 : 0 ] fa_02_13 = fa_01_12 [ 1 ] + fa_01_13 [ 0 ] + b_04_a [  9 ] ;
   wire [ 1 : 0 ] fa_02_14 = fa_01_13 [ 1 ] + fa_01_14 [ 0 ] + b_04_a [ 10 ] ;
   wire [ 1 : 0 ] fa_02_15 = fa_01_14 [ 1 ] + fa_01_15 [ 0 ] + b_04_a [ 11 ] ;
   wire [ 1 : 0 ] fa_02_16 = fa_01_15 [ 1 ] + fa_01_16 [ 0 ] + b_03_a [ 13 ] ;
   wire [ 1 : 0 ] fa_02_17 = fa_01_16 [ 1 ] +  b_02_a [ 15 ] + b_03_a [ 14 ] ;
   
   assign p [ 3 ] = fa_02_03 [ 0 ] ;

   //
   // Row 3
   //
   wire [ 1 : 0 ] fa_03_04 = fa_02_03 [ 1 ] + fa_02_04 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_03_05 = fa_02_04 [ 1 ] + fa_02_05 [ 0 ] + b_05_a [  0 ] ;
   wire [ 1 : 0 ] fa_03_06 = fa_02_05 [ 1 ] + fa_02_06 [ 0 ] + b_05_a [  1 ] ;
   wire [ 1 : 0 ] fa_03_07 = fa_02_06 [ 1 ] + fa_02_07 [ 0 ] + b_05_a [  2 ] ;
   wire [ 1 : 0 ] fa_03_08 = fa_02_07 [ 1 ] + fa_02_08 [ 0 ] + b_05_a [  3 ] ;
   wire [ 1 : 0 ] fa_03_09 = fa_02_08 [ 1 ] + fa_02_09 [ 0 ] + b_05_a [  4 ] ;
   wire [ 1 : 0 ] fa_03_10 = fa_02_09 [ 1 ] + fa_02_10 [ 0 ] + b_05_a [  5 ] ;
   wire [ 1 : 0 ] fa_03_11 = fa_02_10 [ 1 ] + fa_02_11 [ 0 ] + b_05_a [  6 ] ;
   wire [ 1 : 0 ] fa_03_12 = fa_02_11 [ 1 ] + fa_02_12 [ 0 ] + b_05_a [  7 ] ;
   wire [ 1 : 0 ] fa_03_13 = fa_02_12 [ 1 ] + fa_02_13 [ 0 ] + b_05_a [  8 ] ;
   wire [ 1 : 0 ] fa_03_14 = fa_02_13 [ 1 ] + fa_02_14 [ 0 ] + b_05_a [  9 ] ;
   wire [ 1 : 0 ] fa_03_15 = fa_02_14 [ 1 ] + fa_02_15 [ 0 ] + b_05_a [ 10 ] ;
   wire [ 1 : 0 ] fa_03_16 = fa_02_15 [ 1 ] + fa_02_16 [ 0 ] + b_04_a [ 12 ] ;
   wire [ 1 : 0 ] fa_03_17 = fa_02_16 [ 1 ] + fa_02_17 [ 0 ] + b_04_a [ 13 ] ;
   wire [ 1 : 0 ] fa_03_18 = fa_02_17 [ 1 ] +  b_03_a [ 15 ] + b_04_a [ 14 ] ;

   assign p [ 4 ] = fa_03_04 [ 0 ] ;

   //
   // Row 4
   //
   wire [ 1 : 0 ] fa_04_05 = fa_03_04 [ 1 ] + fa_03_05 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_04_06 = fa_03_05 [ 1 ] + fa_03_06 [ 0 ] + b_06_a [  0 ] ;
   wire [ 1 : 0 ] fa_04_07 = fa_03_06 [ 1 ] + fa_03_07 [ 0 ] + b_06_a [  1 ] ;
   wire [ 1 : 0 ] fa_04_08 = fa_03_07 [ 1 ] + fa_03_08 [ 0 ] + b_06_a [  2 ] ;
   wire [ 1 : 0 ] fa_04_09 = fa_03_08 [ 1 ] + fa_03_09 [ 0 ] + b_06_a [  3 ] ;
   wire [ 1 : 0 ] fa_04_10 = fa_03_09 [ 1 ] + fa_03_10 [ 0 ] + b_06_a [  4 ] ;
   wire [ 1 : 0 ] fa_04_11 = fa_03_10 [ 1 ] + fa_03_11 [ 0 ] + b_06_a [  5 ] ;
   wire [ 1 : 0 ] fa_04_12 = fa_03_11 [ 1 ] + fa_03_12 [ 0 ] + b_06_a [  6 ] ;
   wire [ 1 : 0 ] fa_04_13 = fa_03_12 [ 1 ] + fa_03_13 [ 0 ] + b_06_a [  7 ] ;
   wire [ 1 : 0 ] fa_04_14 = fa_03_13 [ 1 ] + fa_03_14 [ 0 ] + b_06_a [  8 ] ;
   wire [ 1 : 0 ] fa_04_15 = fa_03_14 [ 1 ] + fa_03_15 [ 0 ] + b_06_a [  9 ] ;
   wire [ 1 : 0 ] fa_04_16 = fa_03_15 [ 1 ] + fa_03_16 [ 0 ] + b_05_a [ 11 ] ;
   wire [ 1 : 0 ] fa_04_17 = fa_03_16 [ 1 ] + fa_03_17 [ 0 ] + b_05_a [ 12 ] ;
   wire [ 1 : 0 ] fa_04_18 = fa_03_17 [ 1 ] + fa_03_18 [ 0 ] + b_05_a [ 13 ] ;
   wire [ 1 : 0 ] fa_04_19 = fa_03_18 [ 1 ] +  b_04_a [ 15 ] + b_05_a [ 14 ] ;

    assign p [ 5 ] = fa_04_05 [ 0 ] ;


   //
   // Row 5
   //
   wire [ 1 : 0 ] fa_05_06 = fa_04_05 [ 1 ] + fa_04_06 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_05_07 = fa_04_06 [ 1 ] + fa_04_07 [ 0 ] + b_07_a [  0 ] ;
   wire [ 1 : 0 ] fa_05_08 = fa_04_07 [ 1 ] + fa_04_08 [ 0 ] + b_07_a [  1 ] ;
   wire [ 1 : 0 ] fa_05_09 = fa_04_08 [ 1 ] + fa_04_09 [ 0 ] + b_07_a [  2 ] ;
   wire [ 1 : 0 ] fa_05_10 = fa_04_09 [ 1 ] + fa_04_10 [ 0 ] + b_07_a [  3 ] ;
   wire [ 1 : 0 ] fa_05_11 = fa_04_10 [ 1 ] + fa_04_11 [ 0 ] + b_07_a [  4 ] ;
   wire [ 1 : 0 ] fa_05_12 = fa_04_11 [ 1 ] + fa_04_12 [ 0 ] + b_07_a [  5 ] ;
   wire [ 1 : 0 ] fa_05_13 = fa_04_12 [ 1 ] + fa_04_13 [ 0 ] + b_07_a [  6 ] ;
   wire [ 1 : 0 ] fa_05_14 = fa_04_13 [ 1 ] + fa_04_14 [ 0 ] + b_07_a [  7 ] ;
   wire [ 1 : 0 ] fa_05_15 = fa_04_14 [ 1 ] + fa_04_15 [ 0 ] + b_07_a [  8 ] ;
   wire [ 1 : 0 ] fa_05_16 = fa_04_15 [ 1 ] + fa_04_16 [ 0 ] + b_06_a [ 10 ] ;
   wire [ 1 : 0 ] fa_05_17 = fa_04_16 [ 1 ] + fa_04_17 [ 0 ] + b_06_a [ 11 ] ;
   wire [ 1 : 0 ] fa_05_18 = fa_04_17 [ 1 ] + fa_04_18 [ 0 ] + b_06_a [ 12 ] ;
   wire [ 1 : 0 ] fa_05_19 = fa_04_18 [ 1 ] + fa_04_19 [ 0 ] + b_06_a [ 13 ] ;
   wire [ 1 : 0 ] fa_05_20 = fa_04_19 [ 1 ] +  b_05_a [ 15 ] + b_06_a [ 14 ] ;

   assign p [ 6 ] = fa_05_06 [ 0 ] ;


   //
   // Row 6
   //
   wire [ 1 : 0 ] fa_06_07 = fa_05_06 [ 1 ] + fa_05_07 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_06_08 = fa_05_07 [ 1 ] + fa_05_08 [ 0 ] + b_08_a [  0 ] ;
   wire [ 1 : 0 ] fa_06_09 = fa_05_08 [ 1 ] + fa_05_09 [ 0 ] + b_08_a [  1 ] ;
   wire [ 1 : 0 ] fa_06_10 = fa_05_09 [ 1 ] + fa_05_10 [ 0 ] + b_08_a [  2 ] ;
   wire [ 1 : 0 ] fa_06_11 = fa_05_10 [ 1 ] + fa_05_11 [ 0 ] + b_08_a [  3 ] ;
   wire [ 1 : 0 ] fa_06_12 = fa_05_11 [ 1 ] + fa_05_12 [ 0 ] + b_08_a [  4 ] ;
   wire [ 1 : 0 ] fa_06_13 = fa_05_12 [ 1 ] + fa_05_13 [ 0 ] + b_08_a [  5 ] ;
   wire [ 1 : 0 ] fa_06_14 = fa_05_13 [ 1 ] + fa_05_14 [ 0 ] + b_08_a [  6 ] ;
   wire [ 1 : 0 ] fa_06_15 = fa_05_14 [ 1 ] + fa_05_15 [ 0 ] + b_08_a [  7 ] ;
   wire [ 1 : 0 ] fa_06_16 = fa_05_15 [ 1 ] + fa_05_16 [ 0 ] + b_07_a [  9 ] ;
   wire [ 1 : 0 ] fa_06_17 = fa_05_16 [ 1 ] + fa_05_17 [ 0 ] + b_07_a [ 10 ] ;
   wire [ 1 : 0 ] fa_06_18 = fa_05_17 [ 1 ] + fa_05_18 [ 0 ] + b_07_a [ 11 ] ;
   wire [ 1 : 0 ] fa_06_19 = fa_05_18 [ 1 ] + fa_05_19 [ 0 ] + b_07_a [ 12 ] ;
   wire [ 1 : 0 ] fa_06_20 = fa_05_19 [ 1 ] + fa_05_20 [ 0 ] + b_07_a [ 13 ] ;
   wire [ 1 : 0 ] fa_06_21 = fa_05_20 [ 1 ] +  b_06_a [ 15 ] + b_07_a [ 14 ] ;

   assign p [ 7 ] = fa_06_07 [ 0 ] ;


   //
   // Row 7
   //
   wire [ 1 : 0 ] fa_07_08 = fa_06_07 [ 1 ] + fa_06_08 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_07_09 = fa_06_08 [ 1 ] + fa_06_09 [ 0 ] + b_09_a [  0 ] ;
   wire [ 1 : 0 ] fa_07_10 = fa_06_09 [ 1 ] + fa_06_10 [ 0 ] + b_09_a [  1 ] ;
   wire [ 1 : 0 ] fa_07_11 = fa_06_10 [ 1 ] + fa_06_11 [ 0 ] + b_09_a [  2 ] ;
   wire [ 1 : 0 ] fa_07_12 = fa_06_11 [ 1 ] + fa_06_12 [ 0 ] + b_09_a [  3 ] ;
   wire [ 1 : 0 ] fa_07_13 = fa_06_12 [ 1 ] + fa_06_13 [ 0 ] + b_09_a [  4 ] ;
   wire [ 1 : 0 ] fa_07_14 = fa_06_13 [ 1 ] + fa_06_14 [ 0 ] + b_09_a [  5 ] ;
   wire [ 1 : 0 ] fa_07_15 = fa_06_14 [ 1 ] + fa_06_15 [ 0 ] + b_09_a [  6 ] ;
   wire [ 1 : 0 ] fa_07_16 = fa_06_15 [ 1 ] + fa_06_16 [ 0 ] + b_08_a [  8 ] ;
   wire [ 1 : 0 ] fa_07_17 = fa_06_16 [ 1 ] + fa_06_17 [ 0 ] + b_08_a [  9 ] ;
   wire [ 1 : 0 ] fa_07_18 = fa_06_17 [ 1 ] + fa_06_18 [ 0 ] + b_08_a [ 10 ] ;
   wire [ 1 : 0 ] fa_07_19 = fa_06_18 [ 1 ] + fa_06_19 [ 0 ] + b_08_a [ 11 ] ;
   wire [ 1 : 0 ] fa_07_20 = fa_06_19 [ 1 ] + fa_06_20 [ 0 ] + b_08_a [ 12 ] ;
   wire [ 1 : 0 ] fa_07_21 = fa_06_20 [ 1 ] + fa_06_21 [ 0 ] + b_08_a [ 13 ] ;
   wire [ 1 : 0 ] fa_07_22 = fa_06_21 [ 1 ] +  b_07_a [ 15 ] + b_08_a [ 14 ] ;

    assign p [ 8 ] = fa_07_08 [ 0 ] ;


   //
   // Row 8
   //
   wire [ 1 : 0 ] fa_08_09 = fa_07_08 [ 1 ] + fa_07_09 [ 0 ]                 ;
   wire [ 1 : 0 ] fa_08_10 = fa_07_09 [ 1 ] + fa_07_10 [ 0 ] + b_10_a [  0 ] ;
   wire [ 1 : 0 ] fa_08_11 = fa_07_10 [ 1 ] + fa_07_11 [ 0 ] + b_10_a [  1 ] ;
   wire [ 1 : 0 ] fa_08_12 = fa_07_11 [ 1 ] + fa_07_12 [ 0 ] + b_10_a [  2 ] ;
   wire [ 1 : 0 ] fa_08_13 = fa_07_12 [ 1 ] + fa_07_13 [ 0 ] + b_10_a [  3 ] ;
   wire [ 1 : 0 ] fa_08_14 = fa_07_13 [ 1 ] + fa_07_14 [ 0 ] + b_10_a [  4 ] ;
   wire [ 1 : 0 ] fa_08_15 = fa_07_14 [ 1 ] + fa_07_15 [ 0 ] + b_10_a [  5 ] ;
   wire [ 1 : 0 ] fa_08_16 = fa_07_15 [ 1 ] + fa_07_16 [ 0 ] + b_09_a [  7 ] ;
   wire [ 1 : 0 ] fa_08_17 = fa_07_16 [ 1 ] + fa_07_17 [ 0 ] + b_09_a [  8 ] ;
   wire [ 1 : 0 ] fa_08_18 = fa_07_17 [ 1 ] + fa_07_18 [ 0 ] + b_09_a [  9 ] ;
   wire [ 1 : 0 ] fa_08_19 = fa_07_18 [ 1 ] + fa_07_19 [ 0 ] + b_09_a [ 10 ] ;
   wire [ 1 : 0 ] fa_08_20 = fa_07_19 [ 1 ] + fa_07_20 [ 0 ] + b_09_a [ 11 ] ;
   wire [ 1 : 0 ] fa_08_21 = fa_07_20 [ 1 ] + fa_07_21 [ 0 ] + b_09_a [ 12 ] ;
   wire [ 1 : 0 ] fa_08_22 = fa_07_21 [ 1 ] + fa_07_22 [ 0 ] + b_09_a [ 13 ] ;
   wire [ 1 : 0 ] fa_08_23 = fa_07_22 [ 1 ] +  b_08_a [ 15 ] + b_09_a [ 14 ] ;

    assign p [ 9 ] = fa_08_09 [ 0 ] ;


    //
    // Row 9
    //
    wire [ 1 : 0 ] fa_09_10 = fa_08_09 [ 1 ] + fa_08_10 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_09_11 = fa_08_10 [ 1 ] + fa_08_11 [ 0 ] + b_11_a [  0 ] ;
    wire [ 1 : 0 ] fa_09_12 = fa_08_11 [ 1 ] + fa_08_12 [ 0 ] + b_11_a [  1 ] ;
    wire [ 1 : 0 ] fa_09_13 = fa_08_12 [ 1 ] + fa_08_13 [ 0 ] + b_11_a [  2 ] ;
    wire [ 1 : 0 ] fa_09_14 = fa_08_13 [ 1 ] + fa_08_14 [ 0 ] + b_11_a [  3 ] ;
    wire [ 1 : 0 ] fa_09_15 = fa_08_14 [ 1 ] + fa_08_15 [ 0 ] + b_11_a [  4 ] ;
    wire [ 1 : 0 ] fa_09_16 = fa_08_15 [ 1 ] + fa_08_16 [ 0 ] + b_10_a [  6 ] ;
    wire [ 1 : 0 ] fa_09_17 = fa_08_16 [ 1 ] + fa_08_17 [ 0 ] + b_10_a [  7 ] ;
    wire [ 1 : 0 ] fa_09_18 = fa_08_17 [ 1 ] + fa_08_18 [ 0 ] + b_10_a [  8 ] ;
    wire [ 1 : 0 ] fa_09_19 = fa_08_18 [ 1 ] + fa_08_19 [ 0 ] + b_10_a [  9 ] ;
    wire [ 1 : 0 ] fa_09_20 = fa_08_19 [ 1 ] + fa_08_20 [ 0 ] + b_10_a [ 10 ] ;
    wire [ 1 : 0 ] fa_09_21 = fa_08_20 [ 1 ] + fa_08_21 [ 0 ] + b_10_a [ 11 ] ;
    wire [ 1 : 0 ] fa_09_22 = fa_08_21 [ 1 ] + fa_08_22 [ 0 ] + b_10_a [ 12 ] ;
    wire [ 1 : 0 ] fa_09_23 = fa_08_22 [ 1 ] + fa_08_23 [ 0 ] + b_10_a [ 13 ] ; 
    wire [ 1 : 0 ] fa_09_24 = fa_08_23 [ 1 ] +  b_09_a [ 15 ] + b_10_a [ 14 ] ;

    assign p [ 10 ] = fa_09_10 [ 0 ] ;


    //
    // Row 10
    //
    wire [ 1 : 0 ] fa_10_11 = fa_09_10 [ 1 ] + fa_09_11 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_10_12 = fa_09_11 [ 1 ] + fa_09_12 [ 0 ] + b_12_a [  0 ] ;
    wire [ 1 : 0 ] fa_10_13 = fa_09_12 [ 1 ] + fa_09_13 [ 0 ] + b_12_a [  1 ] ;
    wire [ 1 : 0 ] fa_10_14 = fa_09_13 [ 1 ] + fa_09_14 [ 0 ] + b_12_a [  2 ] ;
    wire [ 1 : 0 ] fa_10_15 = fa_09_14 [ 1 ] + fa_09_15 [ 0 ] + b_12_a [  3 ] ;
    wire [ 1 : 0 ] fa_10_16 = fa_09_15 [ 1 ] + fa_09_16 [ 0 ] + b_11_a [  5 ] ;
    wire [ 1 : 0 ] fa_10_17 = fa_09_16 [ 1 ] + fa_09_17 [ 0 ] + b_11_a [  6 ] ;
    wire [ 1 : 0 ] fa_10_18 = fa_09_17 [ 1 ] + fa_09_18 [ 0 ] + b_11_a [  7 ] ;
    wire [ 1 : 0 ] fa_10_19 = fa_09_18 [ 1 ] + fa_09_19 [ 0 ] + b_11_a [  8 ] ;
    wire [ 1 : 0 ] fa_10_20 = fa_09_19 [ 1 ] + fa_09_20 [ 0 ] + b_11_a [  9 ] ;
    wire [ 1 : 0 ] fa_10_21 = fa_09_20 [ 1 ] + fa_09_21 [ 0 ] + b_11_a [ 10 ] ;
    wire [ 1 : 0 ] fa_10_22 = fa_09_21 [ 1 ] + fa_09_22 [ 0 ] + b_11_a [ 11 ] ;
    wire [ 1 : 0 ] fa_10_23 = fa_09_22 [ 1 ] + fa_09_23 [ 0 ] + b_11_a [ 12 ] ; 
    wire [ 1 : 0 ] fa_10_24 = fa_09_23 [ 1 ] + fa_09_24 [ 0 ] + b_11_a [ 13 ] ;
    wire [ 1 : 0 ] fa_10_25 = fa_09_24 [ 1 ] +  b_10_a [ 15 ] + b_11_a [ 14 ] ;

    assign p [ 11 ] = fa_10_11 [ 0 ] ;

    //
    // Row 11
    //
    wire [ 1 : 0 ] fa_11_12 = fa_10_11 [ 1 ] + fa_10_12 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_11_13 = fa_10_12 [ 1 ] + fa_10_13 [ 0 ] + b_13_a [  0 ] ;
    wire [ 1 : 0 ] fa_11_14 = fa_10_13 [ 1 ] + fa_10_14 [ 0 ] + b_13_a [  1 ] ;
    wire [ 1 : 0 ] fa_11_15 = fa_10_14 [ 1 ] + fa_10_15 [ 0 ] + b_13_a [  2 ] ;
    wire [ 1 : 0 ] fa_11_16 = fa_10_15 [ 1 ] + fa_10_16 [ 0 ] + b_12_a [  4 ] ;
    wire [ 1 : 0 ] fa_11_17 = fa_10_16 [ 1 ] + fa_10_17 [ 0 ] + b_12_a [  5 ] ;
    wire [ 1 : 0 ] fa_11_18 = fa_10_17 [ 1 ] + fa_10_18 [ 0 ] + b_12_a [  6 ] ;
    wire [ 1 : 0 ] fa_11_19 = fa_10_18 [ 1 ] + fa_10_19 [ 0 ] + b_12_a [  7 ] ;
    wire [ 1 : 0 ] fa_11_20 = fa_10_19 [ 1 ] + fa_10_20 [ 0 ] + b_12_a [  8 ] ;
    wire [ 1 : 0 ] fa_11_21 = fa_10_20 [ 1 ] + fa_10_21 [ 0 ] + b_12_a [  9 ] ;
    wire [ 1 : 0 ] fa_11_22 = fa_10_21 [ 1 ] + fa_10_22 [ 0 ] + b_12_a [ 10 ] ;
    wire [ 1 : 0 ] fa_11_23 = fa_10_22 [ 1 ] + fa_10_23 [ 0 ] + b_12_a [ 11 ] ; 
    wire [ 1 : 0 ] fa_11_24 = fa_10_23 [ 1 ] + fa_10_24 [ 0 ] + b_12_a [ 12 ] ;
    wire [ 1 : 0 ] fa_11_25 = fa_10_24 [ 1 ] + fa_10_25 [ 0 ] + b_12_a [ 13 ] ;
    wire [ 1 : 0 ] fa_11_26 = fa_10_25 [ 1 ] +  b_11_a [ 15 ] + b_12_a [ 14 ] ;
    
    assign p [ 12 ] = fa_11_12 [ 0 ] ;

    //
    // Row 12
    //
    wire [ 1 : 0 ] fa_12_13 = fa_11_12 [ 1 ] + fa_11_13 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_12_14 = fa_11_13 [ 1 ] + fa_11_14 [ 0 ] + b_14_a [  0 ] ;
    wire [ 1 : 0 ] fa_12_15 = fa_11_14 [ 1 ] + fa_11_15 [ 0 ] + b_14_a [  1 ] ;
    wire [ 1 : 0 ] fa_12_16 = fa_11_15 [ 1 ] + fa_11_16 [ 0 ] + b_13_a [  3 ] ;
    wire [ 1 : 0 ] fa_12_17 = fa_11_16 [ 1 ] + fa_11_17 [ 0 ] + b_13_a [  4 ] ;
    wire [ 1 : 0 ] fa_12_18 = fa_11_17 [ 1 ] + fa_11_18 [ 0 ] + b_13_a [  5 ] ;
    wire [ 1 : 0 ] fa_12_19 = fa_11_18 [ 1 ] + fa_11_19 [ 0 ] + b_13_a [  6 ] ;
    wire [ 1 : 0 ] fa_12_20 = fa_11_19 [ 1 ] + fa_11_20 [ 0 ] + b_13_a [  7 ] ;
    wire [ 1 : 0 ] fa_12_21 = fa_11_20 [ 1 ] + fa_11_21 [ 0 ] + b_13_a [  8 ] ;
    wire [ 1 : 0 ] fa_12_22 = fa_11_21 [ 1 ] + fa_11_22 [ 0 ] + b_13_a [  9 ] ;
    wire [ 1 : 0 ] fa_12_23 = fa_11_22 [ 1 ] + fa_11_23 [ 0 ] + b_13_a [ 10 ] ; 
    wire [ 1 : 0 ] fa_12_24 = fa_11_23 [ 1 ] + fa_11_24 [ 0 ] + b_13_a [ 11 ] ;
    wire [ 1 : 0 ] fa_12_25 = fa_11_24 [ 1 ] + fa_11_25 [ 0 ] + b_13_a [ 12 ] ;
    wire [ 1 : 0 ] fa_12_26 = fa_11_25 [ 1 ] + fa_11_26 [ 0 ] + b_13_a [ 13 ] ;
    wire [ 1 : 0 ] fa_12_27 = fa_11_26 [ 1 ] +  b_12_a [ 15 ] + b_13_a [ 14 ] ;
    
    assign p [ 13 ] = fa_12_13 [ 0 ] ;

    //
    // Row 13
    //
    wire [ 1 : 0 ] fa_13_14 = fa_12_13 [ 1 ] + fa_12_14 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_13_15 = fa_12_14 [ 1 ] + fa_12_15 [ 0 ] + b_15_a [  0 ] ;
    wire [ 1 : 0 ] fa_13_16 = fa_12_15 [ 1 ] + fa_12_16 [ 0 ] + b_14_a [  2 ] ;
    wire [ 1 : 0 ] fa_13_17 = fa_12_16 [ 1 ] + fa_12_17 [ 0 ] + b_14_a [  3 ] ;
    wire [ 1 : 0 ] fa_13_18 = fa_12_17 [ 1 ] + fa_12_18 [ 0 ] + b_14_a [  4 ] ;
    wire [ 1 : 0 ] fa_13_19 = fa_12_18 [ 1 ] + fa_12_19 [ 0 ] + b_14_a [  5 ] ;
    wire [ 1 : 0 ] fa_13_20 = fa_12_19 [ 1 ] + fa_12_20 [ 0 ] + b_14_a [  6 ] ;
    wire [ 1 : 0 ] fa_13_21 = fa_12_20 [ 1 ] + fa_12_21 [ 0 ] + b_14_a [  7 ] ;
    wire [ 1 : 0 ] fa_13_22 = fa_12_21 [ 1 ] + fa_12_22 [ 0 ] + b_14_a [  8 ] ;
    wire [ 1 : 0 ] fa_13_23 = fa_12_22 [ 1 ] + fa_12_23 [ 0 ] + b_14_a [  9 ] ; 
    wire [ 1 : 0 ] fa_13_24 = fa_12_23 [ 1 ] + fa_12_24 [ 0 ] + b_14_a [ 10 ] ;
    wire [ 1 : 0 ] fa_13_25 = fa_12_24 [ 1 ] + fa_12_25 [ 0 ] + b_14_a [ 11 ] ;
    wire [ 1 : 0 ] fa_13_26 = fa_12_25 [ 1 ] + fa_12_26 [ 0 ] + b_14_a [ 12 ] ;
    wire [ 1 : 0 ] fa_13_27 = fa_12_26 [ 1 ] + fa_12_27 [ 0 ] + b_14_a [ 13 ] ;
    wire [ 1 : 0 ] fa_13_28 = fa_12_27 [ 1 ] +  b_13_a [ 15 ] + b_14_a [ 14 ] ;
    
    assign p [ 14 ] = fa_13_14 [ 0 ] ;


    //
    // Row 14
    //
    wire [ 1 : 0 ] fa_14_15 = fa_13_14 [ 1 ] + fa_13_15 [ 0 ]                 ;
    wire [ 1 : 0 ] fa_14_16 = fa_13_15 [ 1 ] + fa_13_16 [ 0 ] + b_15_a [  1 ] ;
    wire [ 1 : 0 ] fa_14_17 = fa_13_16 [ 1 ] + fa_13_17 [ 0 ] + b_15_a [  2 ] ;
    wire [ 1 : 0 ] fa_14_18 = fa_13_17 [ 1 ] + fa_13_18 [ 0 ] + b_15_a [  3 ] ;
    wire [ 1 : 0 ] fa_14_19 = fa_13_18 [ 1 ] + fa_13_19 [ 0 ] + b_15_a [  4 ] ;
    wire [ 1 : 0 ] fa_14_20 = fa_13_19 [ 1 ] + fa_13_20 [ 0 ] + b_15_a [  5 ] ;
    wire [ 1 : 0 ] fa_14_21 = fa_13_20 [ 1 ] + fa_13_21 [ 0 ] + b_15_a [  6 ] ;
    wire [ 1 : 0 ] fa_14_22 = fa_13_21 [ 1 ] + fa_13_22 [ 0 ] + b_15_a [  7 ] ;
    wire [ 1 : 0 ] fa_14_23 = fa_13_22 [ 1 ] + fa_13_23 [ 0 ] + b_15_a [  8 ] ; 
    wire [ 1 : 0 ] fa_14_24 = fa_13_23 [ 1 ] + fa_13_24 [ 0 ] + b_15_a [  9 ] ;
    wire [ 1 : 0 ] fa_14_25 = fa_13_24 [ 1 ] + fa_13_25 [ 0 ] + b_15_a [ 10 ] ;
    wire [ 1 : 0 ] fa_14_26 = fa_13_25 [ 1 ] + fa_13_26 [ 0 ] + b_15_a [ 11 ] ;
    wire [ 1 : 0 ] fa_14_27 = fa_13_26 [ 1 ] + fa_13_27 [ 0 ] + b_15_a [ 12 ] ;
    wire [ 1 : 0 ] fa_14_28 = fa_13_27 [ 1 ] + fa_13_28 [ 0 ] + b_15_a [ 13 ] ;
    wire [ 1 : 0 ] fa_14_29 = fa_13_28 [ 1 ] +  b_14_a [ 15 ] + b_15_a [ 14 ] ;
    
    assign p [ 15 ] = fa_14_15 [ 0 ] ;


    //
    // Row 15
    //
    wire [ 1 : 0 ] fa_15_16 = fa_14_15 [ 1 ] + fa_14_16 [ 0 ]                  ;
    wire [ 1 : 0 ] fa_15_17 = fa_14_16 [ 1 ] + fa_14_17 [ 0 ] + fa_15_16 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_18 = fa_14_17 [ 1 ] + fa_14_18 [ 0 ] + fa_15_17 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_19 = fa_14_18 [ 1 ] + fa_14_19 [ 0 ] + fa_15_18 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_20 = fa_14_19 [ 1 ] + fa_14_20 [ 0 ] + fa_15_19 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_21 = fa_14_20 [ 1 ] + fa_14_21 [ 0 ] + fa_15_20 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_22 = fa_14_21 [ 1 ] + fa_14_22 [ 0 ] + fa_15_21 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_23 = fa_14_22 [ 1 ] + fa_14_23 [ 0 ] + fa_15_22 [ 1 ] ; 
    wire [ 1 : 0 ] fa_15_24 = fa_14_23 [ 1 ] + fa_14_24 [ 0 ] + fa_15_23 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_25 = fa_14_24 [ 1 ] + fa_14_25 [ 0 ] + fa_15_24 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_26 = fa_14_25 [ 1 ] + fa_14_26 [ 0 ] + fa_15_25 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_27 = fa_14_26 [ 1 ] + fa_14_27 [ 0 ] + fa_15_26 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_28 = fa_14_27 [ 1 ] + fa_14_28 [ 0 ] + fa_15_27 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_29 = fa_14_28 [ 1 ] + fa_14_29 [ 0 ] + fa_15_28 [ 1 ] ;
    wire [ 1 : 0 ] fa_15_30 = fa_14_29 [ 1 ] +  b_15_a [ 15 ] + fa_15_29 [ 1 ] ;
    
    assign p [ 16 ] = fa_15_16 [ 0 ] ;
    assign p [ 17 ] = fa_15_17 [ 0 ] ;
    assign p [ 18 ] = fa_15_18 [ 0 ] ;
    assign p [ 19 ] = fa_15_19 [ 0 ] ;
    assign p [ 20 ] = fa_15_20 [ 0 ] ;
    assign p [ 21 ] = fa_15_21 [ 0 ] ;
    assign p [ 22 ] = fa_15_22 [ 0 ] ;
    assign p [ 23 ] = fa_15_23 [ 0 ] ;
    assign p [ 24 ] = fa_15_24 [ 0 ] ;
    assign p [ 25 ] = fa_15_25 [ 0 ] ;
    assign p [ 26 ] = fa_15_26 [ 0 ] ;
    assign p [ 27 ] = fa_15_27 [ 0 ] ;
    assign p [ 28 ] = fa_15_28 [ 0 ] ;
    assign p [ 29 ] = fa_15_29 [ 0 ] ;
    assign p [ 30 ] = fa_15_30 [ 0 ] ;
    assign p [ 31 ] = fa_15_30 [ 1 ] ;


endmodule
